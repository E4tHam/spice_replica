* a simple RC line ckt
Vin 1 0 PWL 0 5.0e-10 2.0 2e-9 2.0 2.5e-9 0
R_1 1 2 100
C_1 2 0 5e-013
R_2 2 3 100
C_2 3 0 5e-013
R_3 3 4 100
C_3 4 0 5e-013
R_4 4 5 100
C_4 5 0 5e-013
R_5 5 6 100
C_5 6 0 5e-013
R_6 6 7 100
C_6 7 0 5e-013
R_7 7 8 100
C_7 8 0 5e-013
R_8 8 9 100
C_8 9 0 5e-013
R_9 9 10 100
C_9 10 0 5e-013
R_10 10 11 100
C_10 11 0 5e-013
R_11 11 12 100
C_11 12 0 5e-013
R_12 12 13 100
C_12 13 0 5e-013
R_13 13 14 100
C_13 14 0 5e-013
R_14 14 15 100
C_14 15 0 5e-013
R_15 15 16 100
C_15 16 0 5e-013
R_16 16 17 100
C_16 17 0 5e-013
R_17 17 18 100
C_17 18 0 5e-013
R_18 18 19 100
C_18 19 0 5e-013
R_19 19 20 100
C_19 20 0 5e-013
.TRAN TR 1.0e-11 3e-9
.PLOTNV 2
.PLOTNV 10
.PLOTNV 20
.end
