
R1  1 0 1
R2  2 1 1
IDD 0 2 DC 1

.TRAN TR 1 1
.PLOTNV 1 2
