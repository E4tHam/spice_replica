* a RC mesh circuits with two voltage inputs 
Vin1 1 0 PWL 0 3.0e-10 2.0 2e-9 2.0 2.3e-9 0 
Vin2 380 0 PWL 0 8.0e-10 2.0 2.5e-9 2.0 2.8e-9 0 
I0 0 1 dc -0.00185414
R0 1 2 23.7475
I1 0 2 dc -0.00148186
R1 2 3 26.7616
I2 0 3 dc -0.00388652
R2 3 4 24.645
I3 0 4 dc -0.00446097
R3 4 5 14.2192
I4 0 5 dc -0.00536952
R4 5 6 23.6274
I5 0 6 dc -0.00323023
R5 6 7 13.8432
I6 0 7 dc -0.0046626
R6 7 8 11.5056
I7 0 8 dc -0.00297147
R7 8 9 24.4197
I8 0 9 dc -0.00522518
R8 9 10 19.3947
I9 0 10 dc -0.00457769
R9 10 11 7.07511
I10 0 11 dc -0.00327913
R10 11 12 7.74867
I11 0 12 dc -0.00372614
R11 12 13 14.7672
I12 0 13 dc -0.00384293
R12 13 14 28.9767
I13 0 14 dc -0.0053386
R13 14 15 9.07974
I14 0 15 dc -0.00237754
R14 15 16 11.509
I15 0 16 dc -0.00562047
R15 16 17 15.8981
I16 0 17 dc -0.0049473
R16 17 18 8.19043
I17 0 18 dc -0.00141103
R17 18 19 28.5161
I18 0 19 dc -0.00112787
R18 19 20 8.85527
I19 0 21 dc -0.00291091
R19 21 22 8.86842
I20 0 22 dc -0.00364667
R20 22 23 26.9212
I21 0 23 dc -0.00315306
R21 23 24 11.5977
I22 0 24 dc -0.00256797
R22 24 25 24.2523
I23 0 25 dc -0.00153695
R23 25 26 24.2761
I24 0 26 dc -0.00452598
R24 26 27 10.466
I25 0 27 dc -0.00480897
R25 27 28 15.2928
I26 0 28 dc -0.00424413
R26 28 29 28.2489
I27 0 29 dc -0.00351209
R27 29 30 22.186
I28 0 30 dc -0.00318045
R28 30 31 20.2075
I29 0 31 dc -0.00388279
R29 31 32 20.8155
I30 0 32 dc -0.00331713
R30 32 33 20.8061
I31 0 33 dc -0.00169147
R31 33 34 29.019
I32 0 34 dc -0.00172188
R32 34 35 16.1671
I33 0 35 dc -0.00262292
R33 35 36 28.8146
I34 0 36 dc -0.00279092
R34 36 37 14.9552
I35 0 37 dc -0.00150641
R35 37 38 28.8771
I36 0 38 dc -0.00592308
R36 38 39 19.3993
I37 0 39 dc -0.00532957
R37 39 40 8.7469
I38 0 41 dc -0.00554575
R38 41 42 21.2813
I39 0 42 dc -0.0013193
R39 42 43 28.875
I40 0 43 dc -0.00583131
R40 43 44 24.6386
I41 0 44 dc -0.00502582
R41 44 45 19.2813
I42 0 45 dc -0.00241293
R42 45 46 29.0638
I43 0 46 dc -0.00389739
R43 46 47 15.9215
I44 0 47 dc -0.00287718
R44 47 48 28.0852
I45 0 48 dc -0.0011435
R45 48 49 24.2215
I46 0 49 dc -0.00461553
R46 49 50 19.7742
I47 0 50 dc -0.00312944
R47 50 51 21.0536
I48 0 51 dc -0.00473381
R48 51 52 6.72546
I49 0 52 dc -0.00126647
R49 52 53 24.3578
I50 0 53 dc -0.00451752
R50 53 54 8.03166
I51 0 54 dc -0.00251718
R51 54 55 6.8627
I52 0 55 dc -0.0044393
R52 55 56 14.1239
I53 0 56 dc -0.00464722
R53 56 57 9.86465
I54 0 57 dc -0.00177296
R54 57 58 9.04481
I55 0 58 dc -0.00516116
R55 58 59 18.7734
I56 0 59 dc -0.00258572
R56 59 60 18.1934
I57 0 61 dc -0.00316611
R57 61 62 10.342
I58 0 62 dc -0.00464802
R58 62 63 5.03423
I59 0 63 dc -0.00393102
R59 63 64 16.9359
I60 0 64 dc -0.00569929
R60 64 65 24.054
I61 0 65 dc -0.00163867
R61 65 66 5.36946
I62 0 66 dc -0.00349997
R62 66 67 26.1193
I63 0 67 dc -0.00526074
R63 67 68 7.27521
I64 0 68 dc -0.00528876
R64 68 69 24.7234
I65 0 69 dc -0.00389238
R65 69 70 7.48723
I66 0 70 dc -0.00514084
R66 70 71 23.6799
I67 0 71 dc -0.00554186
R67 71 72 17.8036
I68 0 72 dc -0.00542283
R68 72 73 29.0487
I69 0 73 dc -0.00383255
R69 73 74 16.8473
I70 0 74 dc -0.00308778
R70 74 75 21.2586
I71 0 75 dc -0.00540101
R71 75 76 19.6484
I72 0 76 dc -0.00211256
R72 76 77 29.9837
I73 0 77 dc -0.0017959
R73 77 78 22.3899
I74 0 78 dc -0.00450765
R74 78 79 29.6551
I75 0 79 dc -0.00424299
R75 79 80 21.372
I76 0 81 dc -0.00522102
R76 81 82 22.0442
I77 0 82 dc -0.00585074
R77 82 83 13.2915
I78 0 83 dc -0.00500041
R78 83 84 8.98411
I79 0 84 dc -0.0053164
R79 84 85 20.0689
I80 0 85 dc -0.00309979
R80 85 86 29.5339
I81 0 86 dc -0.00534448
R81 86 87 16.6009
I82 0 87 dc -0.00223422
R82 87 88 26.116
I83 0 88 dc -0.00521621
R83 88 89 23.4127
I84 0 89 dc -0.00166097
R84 89 90 16.9201
I85 0 90 dc -0.00492168
R85 90 91 17.4398
I86 0 91 dc -0.00384409
R86 91 92 16.1015
I87 0 92 dc -0.00117614
R87 92 93 13.2962
I88 0 93 dc -0.00313315
R88 93 94 19.5643
I89 0 94 dc -0.00144031
R89 94 95 21.8722
I90 0 95 dc -0.00393718
R90 95 96 10.8927
I91 0 96 dc -0.00472323
R91 96 97 28.9588
I92 0 97 dc -0.00532128
R92 97 98 6.86075
I93 0 98 dc -0.00369905
R93 98 99 14.5704
I94 0 99 dc -0.00100923
R94 99 100 22.9154
I95 0 101 dc -0.00126829
R95 101 102 5.52612
I96 0 102 dc -0.00479281
R96 102 103 20.724
I97 0 103 dc -0.00565507
R97 103 104 18.6985
I98 0 104 dc -0.00307017
R98 104 105 14.824
I99 0 105 dc -0.0019879
R99 105 106 12.7021
I100 0 106 dc -0.00204625
R100 106 107 20.2773
I101 0 107 dc -0.0028597
R101 107 108 9.01626
I102 0 108 dc -0.00330112
R102 108 109 25.0745
I103 0 109 dc -0.00191713
R103 109 110 22.9484
I104 0 110 dc -0.00338343
R104 110 111 8.54386
I105 0 111 dc -0.00416829
R105 111 112 11.0641
I106 0 112 dc -0.00162075
R106 112 113 26.787
I107 0 113 dc -0.00151705
R107 113 114 23.8602
I108 0 114 dc -0.0029029
R108 114 115 18.9184
I109 0 115 dc -0.00139119
R109 115 116 14.4344
I110 0 116 dc -0.00412592
R110 116 117 24.7405
I111 0 117 dc -0.0031068
R111 117 118 25.6061
I112 0 118 dc -0.00375958
R112 118 119 23.205
I113 0 119 dc -0.00344407
R113 119 120 11.5546
I114 0 121 dc -0.00348955
R114 121 122 17.2392
I115 0 122 dc -0.00345751
R115 122 123 26.2393
I116 0 123 dc -0.00559449
R116 123 124 14.049
I117 0 124 dc -0.00372895
R117 124 125 20.1133
I118 0 125 dc -0.00404829
R118 125 126 16.0205
I119 0 126 dc -0.00453361
R119 126 127 10.4038
I120 0 127 dc -0.0048284
R120 127 128 12.6597
I121 0 128 dc -0.00493122
R121 128 129 7.24479
I122 0 129 dc -0.00549298
R122 129 130 28.3397
I123 0 130 dc -0.00583691
R123 130 131 20.4637
I124 0 131 dc -0.0013346
R124 131 132 7.82577
I125 0 132 dc -0.00415328
R125 132 133 6.85538
I126 0 133 dc -0.00378704
R126 133 134 10.8551
I127 0 134 dc -0.00405981
R127 134 135 28.3638
I128 0 135 dc -0.00385851
R128 135 136 19.3565
I129 0 136 dc -0.00332216
R129 136 137 8.02135
I130 0 137 dc -0.00218092
R130 137 138 29.9652
I131 0 138 dc -0.0037861
R131 138 139 26.5945
I132 0 139 dc -0.0024356
R132 139 140 23.2486
I133 0 141 dc -0.00510629
R133 141 142 17.2183
I134 0 142 dc -0.00396524
R134 142 143 7.80402
I135 0 143 dc -0.0017915
R135 143 144 22.4767
I136 0 144 dc -0.00397411
R136 144 145 27.0748
I137 0 145 dc -0.00315551
R137 145 146 10.252
I138 0 146 dc -0.00191088
R138 146 147 22.1871
I139 0 147 dc -0.00209063
R139 147 148 11.6116
I140 0 148 dc -0.0021155
R140 148 149 17.3164
I141 0 149 dc -0.00233909
R141 149 150 16.1514
I142 0 150 dc -0.00218124
R142 150 151 12.4197
I143 0 151 dc -0.00425315
R143 151 152 23.7441
I144 0 152 dc -0.00446295
R144 152 153 15.6223
I145 0 153 dc -0.00479778
R145 153 154 14.9599
I146 0 154 dc -0.00286996
R146 154 155 21.0274
I147 0 155 dc -0.00366909
R147 155 156 27.4797
I148 0 156 dc -0.00427696
R148 156 157 28.2667
I149 0 157 dc -0.00104914
R149 157 158 9.31118
I150 0 158 dc -0.00421691
R150 158 159 24.151
I151 0 159 dc -0.00438168
R151 159 160 24.2622
I152 0 161 dc -0.0047774
R152 161 162 27.3984
I153 0 162 dc -0.00208905
R153 162 163 20.915
I154 0 163 dc -0.00398595
R154 163 164 20.558
I155 0 164 dc -0.00282598
R155 164 165 6.77297
I156 0 165 dc -0.00226244
R156 165 166 14.0275
I157 0 166 dc -0.00341815
R157 166 167 17.5926
I158 0 167 dc -0.00244955
R158 167 168 10.9678
I159 0 168 dc -0.00431243
R159 168 169 27.4424
I160 0 169 dc -0.00435725
R160 169 170 6.07954
I161 0 170 dc -0.00518805
R161 170 171 19.3007
I162 0 171 dc -0.00191918
R162 171 172 5.661
I163 0 172 dc -0.00337658
R163 172 173 19.0792
I164 0 173 dc -0.00183949
R164 173 174 20.261
I165 0 174 dc -0.00421055
R165 174 175 12.6598
I166 0 175 dc -0.00578392
R166 175 176 24.1488
I167 0 176 dc -0.00417999
R167 176 177 6.71749
I168 0 177 dc -0.00165327
R168 177 178 23.9281
I169 0 178 dc -0.00340159
R169 178 179 22.8674
I170 0 179 dc -0.00157633
R170 179 180 21.0167
I171 0 181 dc -0.00299175
R171 181 182 22.6573
I172 0 182 dc -0.00491981
R172 182 183 22.6266
I173 0 183 dc -0.0023427
R173 183 184 24.5119
I174 0 184 dc -0.00167071
R174 184 185 11.923
I175 0 185 dc -0.00140627
R175 185 186 10.3315
I176 0 186 dc -0.00198045
R176 186 187 20.4802
I177 0 187 dc -0.00403361
R177 187 188 18.7327
I178 0 188 dc -0.00383768
R178 188 189 8.13408
I179 0 189 dc -0.00136006
R179 189 190 27.0709
I180 0 190 dc -0.00176638
R180 190 191 19.1444
I181 0 191 dc -0.00258311
R181 191 192 13.3699
I182 0 192 dc -0.00202796
R182 192 193 21.9067
I183 0 193 dc -0.00119869
R183 193 194 6.05931
I184 0 194 dc -0.00507981
R184 194 195 6.61576
I185 0 195 dc -0.00453901
R185 195 196 15.2378
I186 0 196 dc -0.00543924
R186 196 197 28.492
I187 0 197 dc -0.00101511
R187 197 198 13.7694
I188 0 198 dc -0.00569214
R188 198 199 29.7856
I189 0 199 dc -0.00279359
R189 199 200 29.4184
I190 0 201 dc -0.00113172
R190 201 202 13.5272
I191 0 202 dc -0.00523098
R191 202 203 15.9554
I192 0 203 dc -0.0045176
R192 203 204 19.2651
I193 0 204 dc -0.00151733
R193 204 205 9.52156
I194 0 205 dc -0.00220111
R194 205 206 22.1062
I195 0 206 dc -0.00592553
R195 206 207 17.8402
I196 0 207 dc -0.00550448
R196 207 208 16.6705
I197 0 208 dc -0.00337179
R197 208 209 15.1883
I198 0 209 dc -0.00479246
R198 209 210 7.87561
I199 0 210 dc -0.00172933
R199 210 211 22.4783
I200 0 211 dc -0.00230096
R200 211 212 18.2552
I201 0 212 dc -0.00133151
R201 212 213 8.72045
I202 0 213 dc -0.0030435
R202 213 214 7.08991
I203 0 214 dc -0.00419548
R203 214 215 5.40547
I204 0 215 dc -0.00219926
R204 215 216 19.5024
I205 0 216 dc -0.00180503
R205 216 217 11.6156
I206 0 217 dc -0.00138355
R206 217 218 8.67812
I207 0 218 dc -0.00143658
R207 218 219 8.58887
I208 0 219 dc -0.00333878
R208 219 220 23.0508
I209 0 221 dc -0.00338694
R209 221 222 18.9568
I210 0 222 dc -0.00348179
R210 222 223 7.02212
I211 0 223 dc -0.00247308
R211 223 224 12.3838
I212 0 224 dc -0.00265829
R212 224 225 7.11625
I213 0 225 dc -0.00149568
R213 225 226 10.0606
I214 0 226 dc -0.00153832
R214 226 227 9.32931
I215 0 227 dc -0.00517698
R215 227 228 25.6696
I216 0 228 dc -0.00562679
R216 228 229 18.3929
I217 0 229 dc -0.00335571
R217 229 230 22.5237
I218 0 230 dc -0.00354215
R218 230 231 24.193
I219 0 231 dc -0.00591475
R219 231 232 16.5916
I220 0 232 dc -0.00435422
R220 232 233 27.2708
I221 0 233 dc -0.00526831
R221 233 234 23.8236
I222 0 234 dc -0.00458198
R222 234 235 7.17759
I223 0 235 dc -0.0049943
R223 235 236 14.3637
I224 0 236 dc -0.00328572
R224 236 237 14.0894
I225 0 237 dc -0.00488161
R225 237 238 19.9275
I226 0 238 dc -0.00128893
R226 238 239 8.04011
I227 0 239 dc -0.00380277
R227 239 240 21.406
I228 0 241 dc -0.00131671
R228 241 242 18.0635
I229 0 242 dc -0.00521861
R229 242 243 8.94218
I230 0 243 dc -0.00101488
R230 243 244 27.5046
I231 0 244 dc -0.0020859
R231 244 245 9.67967
I232 0 245 dc -0.00583146
R232 245 246 25.4616
I233 0 246 dc -0.00455063
R233 246 247 19.6983
I234 0 247 dc -0.0044054
R234 247 248 24.3437
I235 0 248 dc -0.00216394
R235 248 249 10.4621
I236 0 249 dc -0.00286378
R236 249 250 25.5972
I237 0 250 dc -0.0018144
R237 250 251 20.3043
I238 0 251 dc -0.00161359
R238 251 252 15.8898
I239 0 252 dc -0.0010054
R239 252 253 17.9615
I240 0 253 dc -0.00330613
R240 253 254 22.2003
I241 0 254 dc -0.00116239
R241 254 255 15.1274
I242 0 255 dc -0.00351912
R242 255 256 11.9963
I243 0 256 dc -0.00598699
R243 256 257 14.1064
I244 0 257 dc -0.00285232
R244 257 258 28.7769
I245 0 258 dc -0.00140875
R245 258 259 20.3637
I246 0 259 dc -0.00496598
R246 259 260 13.9022
I247 0 261 dc -0.00585664
R247 261 262 9.56959
I248 0 262 dc -0.00314891
R248 262 263 24.6359
I249 0 263 dc -0.00158759
R249 263 264 18.344
I250 0 264 dc -0.00221353
R250 264 265 20.4136
I251 0 265 dc -0.00488622
R251 265 266 9.58088
I252 0 266 dc -0.00345157
R252 266 267 28.3657
I253 0 267 dc -0.00257545
R253 267 268 13.9914
I254 0 268 dc -0.00150698
R254 268 269 14.3096
I255 0 269 dc -0.00545151
R255 269 270 27.3725
I256 0 270 dc -0.00593565
R256 270 271 7.67525
I257 0 271 dc -0.00174654
R257 271 272 28.3886
I258 0 272 dc -0.00491686
R258 272 273 26.9034
I259 0 273 dc -0.00230925
R259 273 274 8.15823
I260 0 274 dc -0.00369346
R260 274 275 13.68
I261 0 275 dc -0.00292702
R261 275 276 14.2499
I262 0 276 dc -0.0033712
R262 276 277 23.2479
I263 0 277 dc -0.00565448
R263 277 278 17.3951
I264 0 278 dc -0.00336609
R264 278 279 28.9111
I265 0 279 dc -0.00249405
R265 279 280 16.1956
I266 0 281 dc -0.00511011
R266 281 282 14.5576
I267 0 282 dc -0.00463637
R267 282 283 13.7028
I268 0 283 dc -0.00430394
R268 283 284 26.5503
I269 0 284 dc -0.00432521
R269 284 285 25.1238
I270 0 285 dc -0.00562901
R270 285 286 13.0411
I271 0 286 dc -0.00338625
R271 286 287 19.2216
I272 0 287 dc -0.00312751
R272 287 288 28.6557
I273 0 288 dc -0.00144581
R273 288 289 15.6441
I274 0 289 dc -0.00254528
R274 289 290 22.4853
I275 0 290 dc -0.00276928
R275 290 291 18.3786
I276 0 291 dc -0.00156883
R276 291 292 23.4295
I277 0 292 dc -0.00564448
R277 292 293 8.49302
I278 0 293 dc -0.00572227
R278 293 294 5.61351
I279 0 294 dc -0.00300935
R279 294 295 10.0024
I280 0 295 dc -0.00151397
R280 295 296 5.90455
I281 0 296 dc -0.00303131
R281 296 297 16.087
I282 0 297 dc -0.0044153
R282 297 298 11.4527
I283 0 298 dc -0.00505668
R283 298 299 7.47743
I284 0 299 dc -0.00423846
R284 299 300 17.7751
I285 0 301 dc -0.0034983
R285 301 302 8.88332
I286 0 302 dc -0.00416634
R286 302 303 7.68626
I287 0 303 dc -0.00206834
R287 303 304 27.1595
I288 0 304 dc -0.00592974
R288 304 305 5.48297
I289 0 305 dc -0.00530862
R289 305 306 8.01948
I290 0 306 dc -0.0016671
R290 306 307 19.2458
I291 0 307 dc -0.00165463
R291 307 308 26.5903
I292 0 308 dc -0.0037248
R292 308 309 16.086
I293 0 309 dc -0.00258861
R293 309 310 15.7794
I294 0 310 dc -0.00583462
R294 310 311 25.1982
I295 0 311 dc -0.00460709
R295 311 312 26.1412
I296 0 312 dc -0.00565609
R296 312 313 7.87959
I297 0 313 dc -0.0033261
R297 313 314 14.7954
I298 0 314 dc -0.00289928
R298 314 315 11.3232
I299 0 315 dc -0.00166914
R299 315 316 20.5938
I300 0 316 dc -0.00409503
R300 316 317 17.2219
I301 0 317 dc -0.00358852
R301 317 318 24.5359
I302 0 318 dc -0.00239204
R302 318 319 15.644
I303 0 319 dc -0.0015361
R303 319 320 10.8214
I304 0 321 dc -0.00551015
R304 321 322 19.5212
I305 0 322 dc -0.00506614
R305 322 323 24.5536
I306 0 323 dc -0.00453561
R306 323 324 13.574
I307 0 324 dc -0.00567865
R307 324 325 10.1748
I308 0 325 dc -0.00461546
R308 325 326 25.8837
I309 0 326 dc -0.00271847
R309 326 327 13.1706
I310 0 327 dc -0.00269407
R310 327 328 18.27
I311 0 328 dc -0.00377217
R311 328 329 5.39317
I312 0 329 dc -0.00327487
R312 329 330 17.492
I313 0 330 dc -0.00225618
R313 330 331 17.7632
I314 0 331 dc -0.00221593
R314 331 332 20.2497
I315 0 332 dc -0.0024842
R315 332 333 27.8664
I316 0 333 dc -0.00384972
R316 333 334 12.3858
I317 0 334 dc -0.00342591
R317 334 335 8.57683
I318 0 335 dc -0.00421737
R318 335 336 8.31909
I319 0 336 dc -0.00512335
R319 336 337 17.8518
I320 0 337 dc -0.00302892
R320 337 338 8.9524
I321 0 338 dc -0.00458221
R321 338 339 17.0477
I322 0 339 dc -0.00459587
R322 339 340 26.3831
I323 0 341 dc -0.00518482
R323 341 342 16.8165
I324 0 342 dc -0.00556515
R324 342 343 7.09669
I325 0 343 dc -0.00182877
R325 343 344 21.9378
I326 0 344 dc -0.00483875
R326 344 345 27.7672
I327 0 345 dc -0.00314175
R327 345 346 26.4178
I328 0 346 dc -0.00275548
R328 346 347 21.7595
I329 0 347 dc -0.0020897
R329 347 348 17.1997
I330 0 348 dc -0.00199657
R330 348 349 15.2642
I331 0 349 dc -0.0029258
R331 349 350 26.7632
I332 0 350 dc -0.00295118
R332 350 351 24.1784
I333 0 351 dc -0.00383279
R333 351 352 14.3802
I334 0 352 dc -0.00552872
R334 352 353 26.241
I335 0 353 dc -0.00241671
R335 353 354 26.4952
I336 0 354 dc -0.00585881
R336 354 355 24.045
I337 0 355 dc -0.00180734
R337 355 356 9.54384
I338 0 356 dc -0.00359613
R338 356 357 12.7859
I339 0 357 dc -0.00591758
R339 357 358 22.9386
I340 0 358 dc -0.0039038
R340 358 359 15.5035
I341 0 359 dc -0.00308289
R341 359 360 10.1508
I342 0 361 dc -0.00577605
R342 361 362 27.0602
I343 0 362 dc -0.00103126
R343 362 363 7.01397
I344 0 363 dc -0.00246746
R344 363 364 26.7535
I345 0 364 dc -0.00587859
R345 364 365 21.0611
I346 0 365 dc -0.00310391
R346 365 366 26.7298
I347 0 366 dc -0.00257284
R347 366 367 29.8743
I348 0 367 dc -0.0013798
R348 367 368 11.8779
I349 0 368 dc -0.00515875
R349 368 369 5.85182
I350 0 369 dc -0.00480974
R350 369 370 14.5939
I351 0 370 dc -0.0021543
R351 370 371 6.25397
I352 0 371 dc -0.00265311
R352 371 372 29.3944
I353 0 372 dc -0.00473638
R353 372 373 19.932
I354 0 373 dc -0.00410929
R354 373 374 20.3044
I355 0 374 dc -0.00385948
R355 374 375 13.3306
I356 0 375 dc -0.00407488
R356 375 376 14.949
I357 0 376 dc -0.00467476
R357 376 377 5.52033
I358 0 377 dc -0.00293486
R358 377 378 20.3737
I359 0 378 dc -0.00399125
R359 378 379 28.4981
I360 0 379 dc -0.0049439
R360 379 380 25.5136
I361 0 381 dc -0.00510579
R361 381 382 20.41
I362 0 382 dc -0.00254615
R362 382 383 25.5059
I363 0 383 dc -0.00121712
R363 383 384 9.82264
I364 0 384 dc -0.00392944
R364 384 385 9.42803
I365 0 385 dc -0.00319446
R365 385 386 17.5862
I366 0 386 dc -0.00354858
R366 386 387 16.6554
I367 0 387 dc -0.00256587
R367 387 388 9.11201
I368 0 388 dc -0.00476115
R368 388 389 15.6361
I369 0 389 dc -0.00387031
R369 389 390 26.1862
I370 0 390 dc -0.00496459
R370 390 391 8.11511
I371 0 391 dc -0.00563482
R371 391 392 19.4663
I372 0 392 dc -0.00321595
R372 392 393 21.5046
I373 0 393 dc -0.00211966
R373 393 394 5.99472
I374 0 394 dc -0.00265289
R374 394 395 7.3683
I375 0 395 dc -0.00305576
R375 395 396 21.8988
I376 0 396 dc -0.00365837
R376 396 397 6.68531
I377 0 397 dc -0.00508639
R377 397 398 7.65312
I378 0 398 dc -0.00255122
R378 398 399 27.3985
I379 0 399 dc -0.00173761
R379 399 400 9.11553
R380 1 21 26.0594
R381 2 22 5.58403
R382 3 23 29.8221
R383 4 24 19.0277
R384 5 25 19.6515
R385 6 26 12.6468
R386 7 27 8.27178
R387 8 28 28.8252
R388 9 29 7.45773
R389 10 30 8.13235
R390 11 31 18.4091
R391 12 32 14.7299
R392 13 33 10.4472
R393 14 34 14.8293
R394 15 35 9.89796
R395 16 36 29.0146
R396 17 37 18.5598
R397 18 38 22.7248
R398 19 39 13.3698
R399 20 40 25.6101
R400 21 41 18.4956
R401 22 42 24.3829
R402 23 43 5.91001
R403 24 44 28.4682
R404 25 45 24.4972
R405 26 46 16.3793
R406 27 47 28.1137
R407 28 48 8.15837
R408 29 49 6.50589
R409 30 50 27.3952
R410 31 51 11.4557
R411 32 52 27.4382
R412 33 53 14.4194
R413 34 54 5.40606
R414 35 55 19.4934
R415 36 56 20.1351
R416 37 57 6.57216
R417 38 58 16.4925
R418 39 59 24.5937
R419 40 60 15.7782
R420 41 61 8.61533
R421 42 62 10.1304
R422 43 63 27.924
R423 44 64 23.4294
R424 45 65 11.3069
R425 46 66 12.3085
R426 47 67 8.88977
R427 48 68 29.0405
R428 49 69 26.1057
R429 50 70 9.50302
R430 51 71 21.9182
R431 52 72 13.0948
R432 53 73 9.15751
R433 54 74 24.8371
R434 55 75 21.9076
R435 56 76 22.0087
R436 57 77 11.2145
R437 58 78 10.7544
R438 59 79 22.0666
R439 60 80 12.7508
R440 61 81 14.134
R441 62 82 26.1862
R442 63 83 26.5978
R443 64 84 23.8882
R444 65 85 7.98484
R445 66 86 10.6007
R446 67 87 29.4165
R447 68 88 6.05044
R448 69 89 19.9886
R449 70 90 17.9903
R450 71 91 15.0923
R451 72 92 9.90724
R452 73 93 21.8157
R453 74 94 17.894
R454 75 95 24.539
R455 76 96 16.7168
R456 77 97 11.3514
R457 78 98 8.01514
R458 79 99 20.8249
R459 80 100 20.3978
R460 81 101 18.3676
R461 82 102 8.02356
R462 83 103 11.3098
R463 84 104 5.72751
R464 85 105 14.4488
R465 86 106 11.2938
R466 87 107 20.2138
R467 88 108 5.51762
R468 89 109 5.6078
R469 90 110 11.8227
R470 91 111 28.5788
R471 92 112 23.5875
R472 93 113 17.8113
R473 94 114 11.4698
R474 95 115 29.366
R475 96 116 21.6517
R476 97 117 25.8487
R477 98 118 6.21009
R478 99 119 18.4498
R479 100 120 13.2716
R480 101 121 13.8101
R481 102 122 7.89101
R482 103 123 9.39546
R483 104 124 29.19
R484 105 125 25.7703
R485 106 126 20.3075
R486 107 127 21.8566
R487 108 128 5.34198
R488 109 129 29.9528
R489 110 130 8.39822
R490 111 131 5.97976
R491 112 132 15.814
R492 113 133 23.7113
R493 114 134 24.3124
R494 115 135 20.4788
R495 116 136 5.94922
R496 117 137 9.61642
R497 118 138 6.68184
R498 119 139 14.7246
R499 120 140 19.6467
R500 121 141 29.9641
R501 122 142 28.9772
R502 123 143 8.81717
R503 124 144 25.911
R504 125 145 15.3002
R505 126 146 6.54317
R506 127 147 8.75409
R507 128 148 27.6208
R508 129 149 22.4151
R509 130 150 16.1482
R510 131 151 11.421
R511 132 152 9.82907
R512 133 153 13.5365
R513 134 154 23.3892
R514 135 155 13.6978
R515 136 156 26.2014
R516 137 157 11.6341
R517 138 158 20.4526
R518 139 159 7.84526
R519 140 160 23.2531
R520 141 161 9.31831
R521 142 162 5.81434
R522 143 163 17.9095
R523 144 164 9.16527
R524 145 165 21.4373
R525 146 166 13.885
R526 147 167 16.9041
R527 148 168 18.2294
R528 149 169 29.2718
R529 150 170 27.1787
R530 151 171 12.3172
R531 152 172 25.4793
R532 153 173 13.0192
R533 154 174 8.74254
R534 155 175 22.1816
R535 156 176 23.182
R536 157 177 6.82974
R537 158 178 23.6785
R538 159 179 14.7798
R539 160 180 29.4523
R540 161 181 17.9873
R541 162 182 15.0855
R542 163 183 17.564
R543 164 184 16.966
R544 165 185 24.3492
R545 166 186 26.5233
R546 167 187 23.2031
R547 168 188 25.2361
R548 169 189 18.013
R549 170 190 16.6576
R550 171 191 14.7652
R551 172 192 24.1062
R552 173 193 16.4537
R553 174 194 26.4837
R554 175 195 9.9584
R555 176 196 28.4439
R556 177 197 16.3631
R557 178 198 13.992
R558 179 199 9.43087
R559 180 200 8.68599
R560 181 201 10.8816
R561 182 202 19.2537
R562 183 203 17.3332
R563 184 204 24.123
R564 185 205 14.2714
R565 186 206 25.2483
R566 187 207 23.4274
R567 188 208 23.091
R568 189 209 27.7714
R569 190 210 9.78409
R570 191 211 14.8481
R571 192 212 7.56833
R572 193 213 7.96997
R573 194 214 9.18073
R574 195 215 28.3499
R575 196 216 9.82303
R576 197 217 25.628
R577 198 218 27.9865
R578 199 219 9.27454
R579 200 220 27.4967
R580 201 221 10.2096
R581 202 222 5.51929
R582 203 223 9.11353
R583 204 224 9.90331
R584 205 225 22.1764
R585 206 226 26.9815
R586 207 227 7.10227
R587 208 228 9.91664
R588 209 229 23.2701
R589 210 230 25.9624
R590 211 231 21.7357
R591 212 232 24.9588
R592 213 233 5.93524
R593 214 234 23.371
R594 215 235 17.0197
R595 216 236 25.6195
R596 217 237 23.7846
R597 218 238 23.9246
R598 219 239 11.058
R599 220 240 11.9485
R600 221 241 14.616
R601 222 242 21.8507
R602 223 243 21.6973
R603 224 244 24.5976
R604 225 245 13.1841
R605 226 246 23.1607
R606 227 247 7.21207
R607 228 248 9.62607
R608 229 249 14.3936
R609 230 250 18.847
R610 231 251 18.7912
R611 232 252 21.8499
R612 233 253 16.2072
R613 234 254 19.3978
R614 235 255 14.0889
R615 236 256 29.2605
R616 237 257 19.6809
R617 238 258 26.7641
R618 239 259 5.62229
R619 240 260 5.97478
R620 241 261 23.7119
R621 242 262 10.1447
R622 243 263 13.9373
R623 244 264 13.8378
R624 245 265 21.2879
R625 246 266 26.8531
R626 247 267 10.4272
R627 248 268 29.6699
R628 249 269 24.9781
R629 250 270 5.92052
R630 251 271 14.4869
R631 252 272 29.9546
R632 253 273 16.7511
R633 254 274 19.6829
R634 255 275 5.42657
R635 256 276 29.7587
R636 257 277 8.79515
R637 258 278 6.24723
R638 259 279 8.6666
R639 260 280 29.8789
R640 261 281 10.1761
R641 262 282 22.6794
R642 263 283 23.212
R643 264 284 13.6469
R644 265 285 6.89226
R645 266 286 10.8838
R646 267 287 27.0759
R647 268 288 7.80349
R648 269 289 20.1534
R649 270 290 14.2306
R650 271 291 13.1115
R651 272 292 14.1752
R652 273 293 7.68743
R653 274 294 5.94517
R654 275 295 14.8512
R655 276 296 24.1441
R656 277 297 28.1788
R657 278 298 18.4041
R658 279 299 18.2643
R659 280 300 5.67766
R660 281 301 7.90649
R661 282 302 15.7455
R662 283 303 7.4692
R663 284 304 9.84676
R664 285 305 16.5393
R665 286 306 13.4159
R666 287 307 27.1058
R667 288 308 15.6847
R668 289 309 19.3552
R669 290 310 19.4325
R670 291 311 14.3267
R671 292 312 14.0589
R672 293 313 8.80877
R673 294 314 5.60558
R674 295 315 29.8467
R675 296 316 9.11243
R676 297 317 8.01488
R677 298 318 21.7386
R678 299 319 19.6489
R679 300 320 23.1932
R680 301 321 12.9386
R681 302 322 13.8201
R682 303 323 16.313
R683 304 324 14.9731
R684 305 325 12.6763
R685 306 326 14.4645
R686 307 327 27.389
R687 308 328 7.36617
R688 309 329 26.4261
R689 310 330 6.79327
R690 311 331 11.2098
R691 312 332 9.60675
R692 313 333 20.5261
R693 314 334 19.6331
R694 315 335 10.3028
R695 316 336 16.4275
R696 317 337 20.1973
R697 318 338 28.3173
R698 319 339 6.46745
R699 320 340 15.1888
R700 321 341 17.4574
R701 322 342 16.6014
R702 323 343 23.3116
R703 324 344 27.3172
R704 325 345 22.648
R705 326 346 6.74562
R706 327 347 17.8339
R707 328 348 17.7983
R708 329 349 6.38772
R709 330 350 23.8066
R710 331 351 7.59542
R711 332 352 12.2798
R712 333 353 27.756
R713 334 354 26.6425
R714 335 355 14.2902
R715 336 356 5.64634
R716 337 357 22.5383
R717 338 358 6.23158
R718 339 359 19.602
R719 340 360 28.5486
R720 341 361 26.297
R721 342 362 16.1993
R722 343 363 19.1817
R723 344 364 25.1569
R724 345 365 20.4511
R725 346 366 12.1271
R726 347 367 18.2989
R727 348 368 24.47
R728 349 369 6.97572
R729 350 370 24.3739
R730 351 371 11.1801
R731 352 372 25.4719
R732 353 373 13.5045
R733 354 374 7.00179
R734 355 375 9.5505
R735 356 376 14.6827
R736 357 377 19.7191
R737 358 378 26.5796
R738 359 379 11.3257
R739 360 380 10.6048
R740 361 381 12.8231
R741 362 382 19.4008
R742 363 383 28.4588
R743 364 384 22.8855
R744 365 385 11.4684
R745 366 386 7.14665
R746 367 387 29.4296
R747 368 388 17.9106
R748 369 389 13.7754
R749 370 390 16.5349
R750 371 391 13.8702
R751 372 392 24.9359
R752 373 393 10.5538
R753 374 394 20.7137
R754 375 395 9.06278
R755 376 396 16.7552
R756 377 397 14.697
R757 378 398 13.3912
R758 379 399 19.0221
R759 380 400 22.5033
V1 9 0 dc 1.8
V2 17 0 dc 1.8
V3 161 0 dc 1.8
V4 169 0 dc 1.8
V5 177 0 dc 1.8
V6 321 0 dc 1.8
V7 329 0 dc 1.8
V8 337 0 dc 1.8
C1 6 0 1.40249e-12
C2 11 0 1.21309e-12
C3 16 0 2.30534e-12
C4 101 0 2.42177e-12
C5 106 0 1.61999e-12
C6 111 0 1.42276e-12
C7 116 0 1.72926e-12
C8 201 0 2.43442e-12
C9 206 0 1.566e-12
C10 211 0 2.63232e-12
C11 216 0 2.21551e-12
C12 301 0 2.11576e-12
C13 306 0 1.75427e-12
C14 311 0 1.78246e-12
C15 316 0 2.33387e-12
.TRAN TR 1.0e-11 4e-9
.PLOTNV 2
.PLOTNV 40
.PLOTNV 80
.PLOTNV 150
.PLOTNV 200
.PLOTNV 250
.PLOTNV 300
.PLOTNV 375
.end
