* three input nand gate

VDD 110 0 DC 3
Vin1 102 0 PWL 0 5.0e-10 3.0 0.5e-8 3.0 0.6e-8 0.0 1e-8 0.0 1.1e-8 3.0
Vin2 107 0 DC 3
Vin3 108 0 DC 3
M1 104 102 103 n 10e-6 0.35e-6 2
M2 104 102 110 p 90e-6 0.35e-6 1
M3 103 107 109 n 10e-6 0.35e-6 2
M4 104 107 110 p 90e-6 0.35e-6 1
M5 109 108 0 n 10e-6 0.35e-6 2
M6 104 108 110 p 90e-6 0.35e-6 1
C1 104 0 0.1e-12
.MODEL 1 VT -0.75 MU 5e-2 COX 0.3e-4 LAMBDA 0.05 CJ0 4.0e-14
.MODEL 2 VT 0.83 MU 1.5e-1 COX 0.3e-4 LAMBDA 0.05 CJ0 4.0e-14
.TRAN TR 1.0e-11 2.0e-8
.PRINTNV 102
.PRINTNV 104
.PLOTNV 102
.PLOTNV 104
.PLOTBI M1
.PLOTBI M2
.PLOTBI M4
