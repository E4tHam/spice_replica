
* R1  1 0 1
* L1  2 1 1 0
* C1  0 2 1 1

R1  0 1 1
L1  0 1 1 0
C1  0 1 1 1


* VDD 1 0 DC 1
* R1  2 1 1
* L1  3 2 1 0
* C1  0 3 1 10

.DC
