* circuit described in the handout

VDD 103 0 DC 3
Vin 101 0 PWL 0 5.0e-10 3.0
Rin 101 102 10
M1 104 102 103 p 30e-6 0.35e-6 1
M2 104 102 0 n 10e-6 0.35e-6 2
C1 104 0 0.1e-12
.MODEL 1 VT -0.75 MU 5e-2 COX 0.3e-4 LAMBDA 0.05 CJ0 4.0e-14
.MODEL 2 VT 0.83 MU 1.5e-1 COX 0.3e-4 LAMBDA 0.05 CJ0 4.0e-14
.TRAN TR 1.0e-11 2.0e-8
.PLOTNV 102
.PLOTNV 104
.PLOTBI M1
.PLOTBI M2
