
VDD 2 0 DC 2
R1  2 1 1
R2  0 1 1

.DC
.PRINTNV 1 2

* node 2 should be 2
* node 1 should be 1
