
VDD 1 0 DC 1
R1  2 1 1
L1  3 2 1 10
C1  0 3 1 1

.DC
