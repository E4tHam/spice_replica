
R1 1 0 1
L1 1 0 1 100

.DC
